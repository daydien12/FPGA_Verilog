module up_count
(
	input clk, reset, 
	output[3:0] counter
);
	reg [3:0] counter_up;

// up counter
	always @(posedge clk or posedge reset)
	begin
		if(reset)
			counter_up <= 4'd0;
		else
			if(counter_up >= 4'b1110)
				counter_up <= 4'd0;
			else
				counter_up <= counter_up + 1;
		end 
	assign counter = counter_up;
endmodule